module network4x4 #(parameter packet_size=16,xno=4,yno=4)(
input clk,
input i_reset,
input [packet_size-1:0] i_data,
input i_data_valid,
input i_rd_en,
output [packet_size-1:0] o_DATA
);

wire [packet_size-1:0] wire04_1;// 0 sending 	4 receiving
wire [packet_size-1:0] wire04_2;// 0 receiving 	4 sending
wire [packet_size-1:0] wire01_1;// 0 sending 	1 receiving
wire [packet_size-1:0] wire01_2;// 0 receiving 	1 sending
wire [packet_size-1:0] wire15_1;// 1 sending 	5 receiving
wire [packet_size-1:0] wire15_2;// 1 receiving 	5 sending
wire [packet_size-1:0] wire45_1;// 4 sending	5 receiving
wire [packet_size-1:0] wire45_2;// 4 receiving 	5 sending

wire [packet_size-1:0] wire8C_1;// 8 sending 	C receiving
wire [packet_size-1:0] wire8C_2;// 8 receiving 	C sending
wire [packet_size-1:0] wire89_1;// 8 sending 	9 receiving
wire [packet_size-1:0] wire89_2;// 8 receiving 	9 sending
wire [packet_size-1:0] wire9D_1;// 9 sending 	D receiving
wire [packet_size-1:0] wire9D_2;// 9 receiving 	D sending
wire [packet_size-1:0] wireCD_1;// C sending	D receiving
wire [packet_size-1:0] wireCD_2;// C receiving 	D sending

wire [packet_size-1:0] wire26_1;
wire [packet_size-1:0] wire26_2;
wire [packet_size-1:0] wire23_1;
wire [packet_size-1:0] wire23_2;
wire [packet_size-1:0] wire37_1;
wire [packet_size-1:0] wire37_2;
wire [packet_size-1:0] wire67_1;
wire [packet_size-1:0] wire67_2;

wire [packet_size-1:0] wireAE_1;
wire [packet_size-1:0] wireAE_2;
wire [packet_size-1:0] wireAB_1;
wire [packet_size-1:0] wireAB_2;
wire [packet_size-1:0] wireBF_1;
wire [packet_size-1:0] wireBF_2;
wire [packet_size-1:0] wireEF_1;
wire [packet_size-1:0] wireEF_2;

wire [packet_size-1:0] wire12_1;
wire [packet_size-1:0] wire12_2;
wire [packet_size-1:0] wire56_1;
wire [packet_size-1:0] wire56_2;
wire [packet_size-1:0] wire9A_1;
wire [packet_size-1:0] wire9A_2;
wire [packet_size-1:0] wireDE_1;
wire [packet_size-1:0] wireDE_2;

wire [packet_size-1:0] wire48_1;
wire [packet_size-1:0] wire48_2;
wire [packet_size-1:0] wire59_1;
wire [packet_size-1:0] wire59_2;
wire [packet_size-1:0] wire6A_1;
wire [packet_size-1:0] wire6A_2;
wire [packet_size-1:0] wire7B_1;
wire [packet_size-1:0] wire7B_2;

wire [48:0] data_valid;
wire [48:0] ready;

switch #(.packet_size(16),.x(2'd0),.y(2'd0), .RTfile("RTinitialize.h"), .numWeight(10)) switch0(
.clk(clk),
.i_data_left(i_data),//dataIn_left
.i_data_right(wire04_2), //dataIn_right
.i_data_up(wire01_2),
.i_data_down(),
.i_wr_valid_left(i_data_valid),
.i_wr_valid_right(data_valid[7]),
.i_wr_valid_up(data_valid[1]),
.i_wr_valid_down(1'b0),
.i_reset(i_reset), // Assigning a single reset signal for the entire circuit, to be kept high for sometime for circuit initialization
.o_data_left(), //dataOut_left
.o_data_right(wire04_1),
.o_data_up(wire01_1),
.o_data_down(),
.i_rd_fifoReady_left(1'b0), // given by an external module
.i_rd_fifoReady_right(ready[7]),
.i_rd_fifoReady_up(ready[1]),
.i_rd_fifoReady_down(1'b0),
.o_rd_valid_left(), //data_valid_left
.o_rd_valid_right(data_valid[6]), //data_valid_right
.o_rd_valid_up(data_valid[0]),
.o_rd_valid_down(),

.o_wr_fifoReady_left(),
.o_wr_fifoReady_right(ready[6]),
.o_wr_fifoReady_up(ready[0]),
.o_wr_fifoReady_down()
);

switch #(.packet_size(16),.x(2'd0),.y(2'd1), .RTfile("rt1.h"), .numWeight(10)) switch1(
.clk(clk),
.i_data_left(),//
.i_data_right(wire15_2),
.i_data_up(wire12_2),//
.i_data_down(wire01_1),

.i_wr_valid_left(1'b0),
.i_wr_valid_right(data_valid[9]),
.i_wr_valid_up(data_valid[3]),
.i_wr_valid_down(data_valid[0]),

.i_reset(i_reset), // Assigning a single reset signal for the entire circuit, to be kept high for sometime for circuit initialization
.o_data_left(), //
.o_data_right(wire15_1),
.o_data_up(wire12_1), // 
.o_data_down(wire01_2),

.i_rd_fifoReady_left(1'b0), // given by an external module
.i_rd_fifoReady_right(ready[9]),
.i_rd_fifoReady_up(ready[3]),
.i_rd_fifoReady_down(ready[0]),

.o_rd_valid_left(),//
.o_rd_valid_right(data_valid[8]),
.o_rd_valid_up(data_valid[2]),
.o_rd_valid_down(data_valid[1]),


.o_wr_fifoReady_left(), //
.o_wr_fifoReady_right(ready[8]), 
.o_wr_fifoReady_up(ready[2]),
.o_wr_fifoReady_down(ready[1])


);

switch #(.packet_size(16),.x(2'd1),.y(2'd0), .RTfile("rt4.h"), .numWeight(10)) switch4(
.clk(clk),
.i_data_left(wire04_1),//dataIn_left
.i_data_right(wire48_2), //dataIn_right 
.i_data_up(wire45_2),
.i_data_down(),//

.i_wr_valid_left(data_valid[6]),
.i_wr_valid_right(data_valid[21]),
.i_wr_valid_up(data_valid[15]),
.i_wr_valid_down(1'b0),

.i_reset(i_reset), // Assigning a single reset signal for the entire circuit, to be kept high for sometime for circuit initialization
.o_data_left(wire04_2), //dataOut_left
.o_data_right(wire48_1),
.o_data_up(wire45_1),
.o_data_down(), // 

.i_rd_fifoReady_left(ready[6]), // given by an external module
.i_rd_fifoReady_right(ready[21]),
.i_rd_fifoReady_up(ready[15]),
.i_rd_fifoReady_down(1'b0),

.o_rd_valid_left(data_valid[7]), //data_valid_left
.o_rd_valid_right(data_valid[20]), //data_valid_right
.o_rd_valid_up(data_valid[14]),
.o_rd_valid_down(), // 


.o_wr_fifoReady_left(ready[7]),
.o_wr_fifoReady_right(ready[20]),
.o_wr_fifoReady_up(ready[14]),
.o_wr_fifoReady_down()


);

switch #(.packet_size(16),.x(2'd1),.y(2'd1), .RTfile("rt5.h"), .numWeight(4)) switch5(
.clk(clk),
.i_data_left(wire15_1),//dataIn_left
.i_data_right(wire59_2), //dataIn_right
.i_data_up(wire56_2),
.i_data_down(wire45_1),//

.i_wr_valid_left(data_valid[8]),
.i_wr_valid_right(data_valid[23]),
.i_wr_valid_up(data_valid[17]),
.i_wr_valid_down(data_valid[14]),

.i_reset(i_reset), // Assigning a single reset signal for the entire circuit, to be kept high for sometime for circuit initialization
.o_data_left(wire15_2), //dataOut_left
.o_data_right(wire59_1),
.o_data_up(wire56_1),
.o_data_down(wire45_2), // 

.i_rd_fifoReady_left(ready[8]), // given by an external module
.i_rd_fifoReady_right(ready[23]),
.i_rd_fifoReady_up(ready[17]),
.i_rd_fifoReady_down(ready[14]),

.o_rd_valid_left(data_valid[9]), //data_valid_left
.o_rd_valid_right(data_valid[22]), //data_valid_right
.o_rd_valid_up(data_valid[16]),
.o_rd_valid_down(data_valid[15]), // 


.o_wr_fifoReady_left(ready[9]),
.o_wr_fifoReady_right(ready[22]),
.o_wr_fifoReady_up(ready[16]),
.o_wr_fifoReady_down(ready[15])


);

switch #(.packet_size(16),.x(2'd2),.y(2'd0), .RTfile("rt8.h"), .numWeight(3)) switch8(
.clk(clk),
.i_data_left(wire48_1),
.i_data_right(wire8C_2), //
.i_data_up(wire89_2),
.i_data_down(),//

.i_wr_valid_left(data_valid[20]),
.i_wr_valid_right(data_valid[35]),
.i_wr_valid_up(data_valid[29]),
.i_wr_valid_down(1'b0),

.i_reset(i_reset), // Assigning a single reset signal for the entire circuit, to be kept high for sometime for circuit initialization
.o_data_left(wire48_2),
.o_data_right(wire8C_1), // 
.o_data_up(wire89_1),
.o_data_down(), // 

.i_rd_fifoReady_left(ready[20]), // given by an external module
.i_rd_fifoReady_right(ready[35]),
.i_rd_fifoReady_up(ready[29]),
.i_rd_fifoReady_down(1'b0),

.o_rd_valid_left(data_valid[21]), //data_valid_left
.o_rd_valid_right(data_valid[34]), //
.o_rd_valid_up(data_valid[28]),
.o_rd_valid_down(), //


.o_wr_fifoReady_left(ready[21]),
.o_wr_fifoReady_right(ready[34]),//
.o_wr_fifoReady_up(ready[28]),
.o_wr_fifoReady_down()


);

switch #(.packet_size(16),.x(2'd2),.y(2'd1), .RTfile("rt9.h"), .numWeight(3)) switch9(

.clk(clk),
.i_data_left(wire59_1),
.i_data_right(wire9D_2),//
.i_data_up(wire9A_2),//
.i_data_down(wire89_1),

.i_wr_valid_left(data_valid[22]),
.i_wr_valid_right(data_valid[37]),
.i_wr_valid_up(data_valid[31]),
.i_wr_valid_down(data_valid[28]),

.i_reset(i_reset), // Assigning a single reset signal for the entire circuit, to be kept high for sometime for circuit initialization
.o_data_left(wire59_2),
.o_data_right(wire9D_1), //
.o_data_up(wire9A_1),//
.o_data_down(wire89_2),

.i_rd_fifoReady_left(ready[22]), // given by an external module
.i_rd_fifoReady_right(ready[37]),
.i_rd_fifoReady_up(ready[31]),
.i_rd_fifoReady_down(ready[28]),

.o_rd_valid_left(data_valid[23]),
.o_rd_valid_right(data_valid[36]), //
.o_rd_valid_up(data_valid[30]),//
.o_rd_valid_down(data_valid[29]),


.o_wr_fifoReady_left(ready[23]),
.o_wr_fifoReady_right(ready[36]),//
.o_wr_fifoReady_up(ready[30]),//
.o_wr_fifoReady_down(ready[29])


);

switch #(.packet_size(16),.x(2'd3),.y(2'd0), .RTfile("rt12.h"), .numWeight(10)) switchC(
.clk(clk),
.i_data_left(wire8C_1),//dataIn_left
.i_data_right(), //dataIn_right
.i_data_up(wireCD_2),
.i_data_down(),//

.i_wr_valid_left(data_valid[34]),
.i_wr_valid_right(1'b0),
.i_wr_valid_up(data_valid[43]),
.i_wr_valid_down(1'b0),

.i_reset(i_reset), // Assigning a single reset signal for the entire circuit, to be kept high for sometime for circuit initialization
.o_data_left(wire8C_2), //dataOut_left
.o_data_right(),
.o_data_up(wireCD_1),
.o_data_down(), // 

.i_rd_fifoReady_left(ready[34]), // given by an external module
.i_rd_fifoReady_right(1'b0),
.i_rd_fifoReady_up(ready[43]),
.i_rd_fifoReady_down(1'b0),

.o_rd_valid_left(data_valid[35]), //data_valid_left
.o_rd_valid_right(), //data_valid_right
.o_rd_valid_up(data_valid[42]),
.o_rd_valid_down(), // 


.o_wr_fifoReady_left(ready[35]),
.o_wr_fifoReady_right(),
.o_wr_fifoReady_up(ready[42]),
.o_wr_fifoReady_down()


);

switch #(.packet_size(16),.x(2'd3),.y(2'd1), .RTfile("rt13.h"), .numWeight(10)) switchD(
.clk(clk),
.i_data_left(wire9D_1),//dataIn_left
.i_data_right(), //dataIn_right
.i_data_up(wireDE_2),
.i_data_down(wireCD_1),

.i_wr_valid_left(data_valid[36]),
.i_wr_valid_right(1'b0),
.i_wr_valid_up(data_valid[45]),
.i_wr_valid_down(data_valid[42]),

.i_reset(i_reset), // Assigning a single reset signal for the entire circuit, to be kept high for sometime for circuit initialization
.o_data_left(wire9D_2), //dataOut_left
.o_data_right(),
.o_data_up(wireDE_1),
.o_data_down(wireCD_2),

.i_rd_fifoReady_left(ready[36]), // given by an external module
.i_rd_fifoReady_right(1'b0),
.i_rd_fifoReady_up(ready[45]),
.i_rd_fifoReady_down(ready[42]),

.o_rd_valid_left(data_valid[37]), //data_valid_left
.o_rd_valid_right(), //data_valid_right
.o_rd_valid_up(data_valid[44]),
.o_rd_valid_down(data_valid[43]),


.o_wr_fifoReady_left(ready[37]),
.o_wr_fifoReady_right(),
.o_wr_fifoReady_up(ready[44]),
.o_wr_fifoReady_down(ready[43])


);

switch #(.packet_size(16),.x(2'd0),.y(2'd2), .RTfile("rt2.h"), .numWeight(10)) switch2(
.clk(clk),
.i_data_left(),//dataIn_left
.i_data_right(wire26_2), //dataIn_right
.i_data_up(wire23_2),
.i_data_down(wire12_1),

.i_wr_valid_left(),
.i_wr_valid_right(data_valid[11]),
.i_wr_valid_up(data_valid[48]),
.i_wr_valid_down(data_valid[2]),

.i_reset(i_reset), // Assigning a single reset signal for the entire circuit, to be kept high for sometime for circuit initialization
.o_data_left(), //dataOut_left
.o_data_right(wire26_1),
.o_data_up(wire23_1),
.o_data_down(wire12_2), // 

.i_rd_fifoReady_left(1'b0), // given by an external module
.i_rd_fifoReady_right(ready[11]),
.i_rd_fifoReady_up(ready[48]),
.i_rd_fifoReady_down(ready[2]),

.o_rd_valid_left(), //data_valid_left
.o_rd_valid_right(data_valid[10]), //data_valid_right
.o_rd_valid_up(data_valid[4]),
.o_rd_valid_down(data_valid[3]), // 


.o_wr_fifoReady_left(),
.o_wr_fifoReady_right(ready[10]),
.o_wr_fifoReady_up(ready[4]),
.o_wr_fifoReady_down(ready[3])


);

switch #(.packet_size(16),.x(2'd0),.y(2'd3), .RTfile("rt3.h"), .numWeight(10)) switch3(
.clk(clk),
.i_data_left(),//dataIn_left
.i_data_right(wire37_2), //dataIn_right
.i_data_up(),
.i_data_down(wire23_1),

.i_wr_valid_left(),
.i_wr_valid_right(data_valid[13]),
.i_wr_valid_up(),
.i_wr_valid_down(data_valid[4]),

.i_reset(i_reset), // Assigning a single reset signal for the entire circuit, to be kept high for sometime for circuit initialization
.o_data_left(), //dataOut_left
.o_data_right(wire37_1),
.o_data_up(),
.o_data_down(wire23_2),

.i_rd_fifoReady_left(1'b0), // given by an external module
.i_rd_fifoReady_right(ready[13]),
.i_rd_fifoReady_up(1'b0),
.i_rd_fifoReady_down(ready[4]),

.o_rd_valid_left(), //data_valid_left
.o_rd_valid_right(data_valid[12]), //data_valid_right
.o_rd_valid_up(),
.o_rd_valid_down(data_valid[48]),


.o_wr_fifoReady_left(),
.o_wr_fifoReady_right(ready[12]),
.o_wr_fifoReady_up(),
.o_wr_fifoReady_down(ready[48])


);

switch #(.packet_size(16),.x(2'd1),.y(2'd2), .RTfile("rt6.h"), .numWeight(4)) switch6(
.clk(clk),
.i_data_left(wire26_1),//dataIn_left
.i_data_right(wire6A_2), //dataIn_right
.i_data_up(wire67_2),
.i_data_down(wire56_1),

.i_wr_valid_left(data_valid[10]),
.i_wr_valid_right(data_valid[25]),
.i_wr_valid_up(data_valid[19]),
.i_wr_valid_down(data_valid[16]),

.i_reset(i_reset), // Assigning a single reset signal for the entire circuit, to be kept high for sometime for circuit initialization
.o_data_left(wire26_2), //dataOut_left
.o_data_right(wire6A_1),
.o_data_up(wire67_1),
.o_data_down(wire56_2),

.i_rd_fifoReady_left(ready[10]), // given by an external module
.i_rd_fifoReady_right(ready[25]),
.i_rd_fifoReady_up(ready[19]),
.i_rd_fifoReady_down(ready[16]),

.o_rd_valid_left(data_valid[11]), //data_valid_left
.o_rd_valid_right(data_valid[24]), //data_valid_right
.o_rd_valid_up(data_valid[18]),
.o_rd_valid_down(data_valid[17]),


.o_wr_fifoReady_left(ready[11]),
.o_wr_fifoReady_right(ready[24]),
.o_wr_fifoReady_up(ready[18]),
.o_wr_fifoReady_down(ready[17])


);

switch #(.packet_size(16),.x(2'd1),.y(2'd3), .RTfile("rt7.h"), .numWeight(4)) switch7(
.clk(clk),
.i_data_left(wire37_1),//dataIn_left
.i_data_right(wire7B_2), //dataIn_right
.i_data_up(),
.i_data_down(wire67_1),

.i_wr_valid_left(data_valid[12]),
.i_wr_valid_right(data_valid[27]),
.i_wr_valid_up(),
.i_wr_valid_down(data_valid[18]),

.i_reset(i_reset), // Assigning a single reset signal for the entire circuit, to be kept high for sometime for circuit initialization
.o_data_left(wire37_2), //dataOut_left
.o_data_right(wire7B_1),
.o_data_up(),
.o_data_down(wire67_2), // 

.i_rd_fifoReady_left(ready[12]), // given by an external module
.i_rd_fifoReady_right(ready[27]),
.i_rd_fifoReady_up(),
.i_rd_fifoReady_down(ready[18]),

.o_rd_valid_left(data_valid[13]), //data_valid_left
.o_rd_valid_right(data_valid[26]), //data_valid_right
.o_rd_valid_up(),
.o_rd_valid_down(data_valid[19]),


.o_wr_fifoReady_left(ready[13]),
.o_wr_fifoReady_right(ready[26]),
.o_wr_fifoReady_up(),
.o_wr_fifoReady_down(ready[19])


);

switch #(.packet_size(16),.x(2'd2),.y(2'd2), .RTfile("rt10.h"), .numWeight(10)) switchA(
.clk(clk),
.i_data_left(wire6A_1),//dataIn_left
.i_data_right(wireAE_2), //dataIn_right
.i_data_up(wireAB_2),
.i_data_down(wire9A_1),

.i_wr_valid_left(data_valid[24]),
.i_wr_valid_right(data_valid[39]),
.i_wr_valid_up(data_valid[33]),
.i_wr_valid_down(data_valid[30]),

.i_reset(i_reset), // Assigning a single reset signal for the entire circuit, to be kept high for sometime for circuit initialization
.o_data_left(wire6A_2), //dataOut_left
.o_data_right(wireAE_1),
.o_data_up(wireAB_1),
.o_data_down(wire9A_2),

.i_rd_fifoReady_left(ready[24]), // given by an external module
.i_rd_fifoReady_right(ready[39]),
.i_rd_fifoReady_up(ready[33]),
.i_rd_fifoReady_down(ready[30]),

.o_rd_valid_left(data_valid[25]), //data_valid_left
.o_rd_valid_right(data_valid[38]), //data_valid_right
.o_rd_valid_up(data_valid[32]),
.o_rd_valid_down(data_valid[31]),


.o_wr_fifoReady_left(ready[25]),
.o_wr_fifoReady_right(ready[38]),
.o_wr_fifoReady_up(ready[32]),
.o_wr_fifoReady_down(ready[31])


);

switch #(.packet_size(16),.x(2'd2),.y(2'd3), .RTfile("rt11.h"), .numWeight(10)) switchB(
.clk(clk),
.i_data_left(wire7B_1),//dataIn_left
.i_data_right(wireBF_2), //dataIn_right
.i_data_up(),
.i_data_down(wireAB_1),

.i_wr_valid_left(data_valid[26]),
.i_wr_valid_right(data_valid[41]),
.i_wr_valid_up(),
.i_wr_valid_down(data_valid[32]),

.i_reset(i_reset), // Assigning a single reset signal for the entire circuit, to be kept high for sometime for circuit initialization
.o_data_left(wire7B_2), //dataOut_left
.o_data_right(wireBF_1),
.o_data_up(),
.o_data_down(wireAB_2),

.i_rd_fifoReady_left(ready[26]), // given by an external module
.i_rd_fifoReady_right(ready[41]),
.i_rd_fifoReady_up(),
.i_rd_fifoReady_down(ready[32]),

.o_rd_valid_left(data_valid[27]), //data_valid_left
.o_rd_valid_right(data_valid[40]), //data_valid_right
.o_rd_valid_up(),
.o_rd_valid_down(data_valid[33]),


.o_wr_fifoReady_left(ready[27]),
.o_wr_fifoReady_right(ready[40]),
.o_wr_fifoReady_up(),
.o_wr_fifoReady_down(ready[33])


);

switch_type_2 #(.packet_size(16),.x(2'd3),.y(2'd2)) switchE(
.clk(clk),
.i_data_left(wireAE_1),//dataIn_left
.i_data_right(), //dataIn_right
.i_data_up(wireEF_2),
.i_data_down(wireDE_1),

.i_wr_valid_left(data_valid[38]),
.i_wr_valid_right(),
.i_wr_valid_up(data_valid[47]),
.i_wr_valid_down(data_valid[44]),

.i_reset(i_reset), // Assigning a single reset signal for the entire circuit, to be kept high for sometime for circuit initialization
.o_data_left(wireAE_2), //dataOut_left
.o_data_right(o_DATA),
.o_data_up(wireEF_1),
.o_data_down(wireDE_2),

.i_rd_fifoReady_left(ready[38]), // given by an external module
.i_rd_fifoReady_right(i_rd_en),
.i_rd_fifoReady_up(ready[47]),
.i_rd_fifoReady_down(ready[44]),

.o_rd_valid_left(data_valid[39]), //data_valid_left
.o_rd_valid_right(), //data_valid_right
.o_rd_valid_up(data_valid[46]),
.o_rd_valid_down(data_valid[45]),


.o_wr_fifoReady_left(ready[39]),
.o_wr_fifoReady_right(),
.o_wr_fifoReady_up(ready[46]),
.o_wr_fifoReady_down(ready[45])

);

switch #(.packet_size(16),.x(2'd3),.y(2'd3), .RTfile("rt15.h"), .numWeight(10)) switchF(
.clk(clk),
.i_data_left(wireBF_1),//dataIn_left
.i_data_right(), //dataIn_right
.i_data_up(),
.i_data_down(wireEF_1),

.i_wr_valid_left(data_valid[40]),
.i_wr_valid_right(),
.i_wr_valid_up(),
.i_wr_valid_down(data_valid[46]),

.i_reset(i_reset), // Assigning a single reset signal for the entire circuit, to be kept high for sometime for circuit initialization
.o_data_left(wireBF_2), //dataOut_left
.o_data_right(),
.o_data_up(),
.o_data_down(wireEF_2),

.i_rd_fifoReady_left(ready[40]), // given by an external module
.i_rd_fifoReady_right(),
.i_rd_fifoReady_up(),
.i_rd_fifoReady_down(ready[46]),

.o_rd_valid_left(data_valid[41]), //data_valid_left
.o_rd_valid_right(), //data_valid_right
.o_rd_valid_up(),
.o_rd_valid_down(data_valid[47]),


.o_wr_fifoReady_left(ready[41]),
.o_wr_fifoReady_right(),
.o_wr_fifoReady_up(),
.o_wr_fifoReady_down(ready[47])


);


endmodule